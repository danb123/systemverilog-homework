//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module halve_tokens
(
    input  clk,
    input  rst,
    input  a,
    output b
);
    // Task:
    // Implement a serial module that reduces amount of incoming '1' tokens by half.
    //
    // Note:
    // Check the waveform diagram in the README for better understanding.
    //
    // Example:
    // a -> 110_011_101_000_1111
    // b -> 010_001_001_000_0101

    logic first_token;

    always_ff @(posedge clk) begin
      if (rst) begin
        first_token <= 0;
      end else if (a && !first_token) begin
        first_token <= 1;
      end else if (b) begin
        first_token <= 0;
      end
    end

    assign b = a && first_token;

endmodule
